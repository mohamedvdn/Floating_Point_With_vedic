library verilog;
use verilog.vl_types.all;
entity M_white_ball is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : out    vl_logic;
        D               : out    vl_logic
    );
end M_white_ball;
